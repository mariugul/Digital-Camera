[aimspice]
[description]
2153
* This is a parametrized testbench for pixel circuit 

.include inc/p18_cmos_models.inc
.include inc/PhotoDiode.inc

.param Ipd_1 	  = 750p 				  ! Photodiode current, range [50 pA, 750 pA]
.param VDD 		  = 1.8 				  ! Supply voltage
.param EXPOSURETIME = 15m 				  ! Exposure time, range [2 ms, 30 ms]

.param TRF        = {EXPOSURETIME/100} 		  ! Risetime and falltime of EXPOSURE and ERASE signals
.param PW         = {EXPOSURETIME} 			  ! Pulsewidth of EXPOSURE and ERASE signals
.param PERIOD     = {EXPOSURETIME*10} 	        ! Period for testbench sources
.param FS = 1k;                   			  ! Sampling clock frequency 
.param CLK_PERIOD = {1/FS} 				  ! Sampling clock period
.param EXPOSE_DLY = {CLK_PERIOD} 			  ! Delay for EXPOSE signalj m
.param NRE_R1_DLY = {2*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE_R1 signal
.param ERASE_DLY  = {6*CLK_PERIOD + EXPOSURETIME} ! Delay for ERASE signal


*TRANSISTORS PARAMETERS - Random values for now
* NMOS Switches 
.param LNswitch = 1.080u
.param WNswitch = 1.080u

* pMOS Switches 
.param LPswitch = 0.36U
.param WPswitch = 1.080U

* Amplifiers 
.param LPamp = 0.36U
.param WPamp = 1.080U

* Active loads 
.param LPload = 0.36U
.param WPload = 1.080U


VDD 1 0 dc VDD
VEXPOSE EXPOSE 0 dc 0 pulse(0 VDD EXPOSE_DLY TRF TRF EXPOSURETIME PERIOD)
VERASE  ERASE  0 dc 0 pulse(0 VDD ERASE_DLY  TRF TRF CLK_PERIOD PERIOD)
VNRE NRE 0 dc 0 pulse(VDD 0 NRE_R1_DLY TRF TRF CLK_PERIOD PERIOD)


************************PIXEL DEFINITION **********************************
*Photodiode
XPD1	1	N1	PhotoDiode	Ipd=750
	
*Expose trigger
M1	N1 	EXPOSE 	N2	0 	NMOS 	L=LNswitch 	W=WNswitch
	
*Erase trigger
M2	N2	ERASE		0	0	NMOS 	L=LNswitch 	W=WNswitch
	
*Sampling Capacitor
Cs	N2	0	2p
	
*Readout circuit
M3 	0 	N2 	N3 	1 	PMOS 	L=LPamp 	W=WPamp
M4 	N3 	NRE	OUT 	1 	PMOS 	L=LPswitch 	W=WPswitch

MC1 	OUT	OUT	1	1 	PMOS 	L=LPload	W=WPload
CC1	OUT	0	3p
****************************************************************************

************************** PLOTS *******************************************
.plot V(N2) V(EXPOSE) V(ERASE)









[dc]
1
VDD
0
1.8
0.1
[tran]
0.01m
60m
0
X
0
[ana]
4 0
[end]
