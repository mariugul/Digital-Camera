//-----------------------------------------------------------------------------
//
// Title       : CTRL_ex_time
// Design      : Digital camera
// Author      : user
// Company     : NTNU
//
//-----------------------------------------------------------------------------
//
// File        : \\sambaad.stud.ntnu.no\mariugul\Documents\Digital_Camera\Digital camera\src\CTRL_ex_time.v
// Generated   : Sat Nov 16 17:13:37 2019
// From        : interface description file
// By          : Itf2Vhdl ver. 1.22
//
//-----------------------------------------------------------------------------
//
// Description : 
//
//-----------------------------------------------------------------------------
`timescale 1 ns / 1 ps

module CTRL_ex_time (Exp_time, Clk, Reset, Exp_increase, Exp_decrease);

output Exp_time;
input Clk, Reset, Exp_increase, Exp_decrease;
wire Clk, Reset, Exp_increase, Exp_decrease, Exp_time;


// -- Enter your statements here -- //		



endmodule
