[aimspice]
[description]
595
*Pixel Circuit 

*<name> <drain> <gate> <source> <bulk> <type> <L>  <W>

.include p18_cmos_models.inc
.include PhotoDiode.inc

.subckt PIXEL VDD VSS EXPOSE ERASE NRE OUT PARAM: Ipd=750p
	* Photodiode
	XPD1	VDD	N1	PhotoDiode	Ipd={Ipd}
	
	*Expose trigger
	MN1 N1 EXPOSE N2 VSS NMOS L=LNswitch W=WNswitch   !Switch 
	*Erase trigger
	MN2 N2 ERASE VSS VSS NMOS L=LNswitch W=WNswitch   !Switch

	*Readout circuit 
	MP3 VSS  N2 N3 1 PMOS L=LPamp W=WPamp     	!Amplifier
	MP4 N3 NRE OUT 1 PMOS L=LPswitch W=WPswitch    	!Switch

	*Sampling capacitor 
	CS N2 VSS 2pf  

.ends PIXEL
[tran]
0.001
0.06
X
X
0
[ana]
4 0
[end]
