//-----------------------------------------------------------------------------
//
// Title       : Timer_counter
// Design      : Digital camera
// Author      : user
// Company     : NTNU
//
//-----------------------------------------------------------------------------
//
// File        : \\sambaad.stud.ntnu.no\mariugul\Documents\Digital_Camera\Digital camera\src\Timer_counter.v
// Generated   : Fri Nov 15 18:49:50 2019
// From        : interface description file
// By          : Itf2Vhdl ver. 1.22
//
//-----------------------------------------------------------------------------
//
// Description : 
//
//-----------------------------------------------------------------------------
`timescale 1 ns / 1 ps

module Timer_counter (Ovf5, Ovf4, Initial, Start, Clk, Reset);

output Ovf5, Ovf4;		   
input Initial, Start, Clk, Reset;
wire Ovf5, Ovf4, Initial, Start, Clk, Reset;

// -- Enter your statements here -- //

endmodule
